module CPU_Top(